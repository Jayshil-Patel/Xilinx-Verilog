`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:34:50 10/06/2020 
// Design Name: 
// Module Name:    swapping_blocking_18ec068 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module swapping_blocking_18ec068(
    );
	 reg[1:0]a;
	 reg[1:0]b;
	 
	 initial begin
	 a=2'b01;
	 b=2'b11;
	 a=a+b;
	 b=a-b;
	 a=a-b;
	 end


endmodule
